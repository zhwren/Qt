/*************************************************************
**                         _ooOoo_                          **
**                        o8888888o                         **
**                        88" . "88                         **
**                        (| -_- |)                         **
**                         O\ = /O                          **
**                     ____/`---'\____                      **
**                   .   ' \\| |// `.                       **
**                    / \\||| : |||// \                     **
**                  / _||||| -:- |||||- \                   **
**                    | | \\\ - /// | |                     **
**                  | \_| ''\---/'' | |                     **
**                   \ .-\__ `-` ___/-. /                   **
**                ___`. .' /--.--\ `. . __                  **
**             ."" '< `.____<|>_/___.' >'"".                **
**            | | : `- \`.;` _ /`;.`/ - ` : | |             **
**              \ \ `-. \_ __\ /__ _/ .-` / /               **
**      ======`-.____`-.___\_____/___.-`____.-'======       **
**                         `=---='                          **
**                                                          **
**      .............................................       **
**             Buddha bless me, No bug forever              **
**                                                          **
**************************************************************
** Author       : generator                                 **
** Email        : zhuhw@ihep.ac.cn/zhwren0211@whu.edu.cn    **
** Last modified: TIME_CONTEXT                       **
** Filename     : demo_xaction.sv
** Discription  :                                           **
*************************************************************/
`ifndef __DEMO_XACTION_SV__
`define __DEMO_XACTION_SV__

`include "demo_dec.sv"
import demo_dec::*;

class demo_xaction extends uvm_sequence_item;
    XACTION_CONTEXT
    extern function new(string name="demo_xaction");
endclass

/*************************************************************
** Time        : TIME_CONTEXT                        **
** Author      : generator                                  **
** Description : Create                                     **
*************************************************************/
function demo_xaction::new(string name="demo_xaction");
    super.new(name);
endfunction

`endif
